#single upper case letter are usually initials
A
B
C
D
E
F
G
H
I
J
K
L
M
N
O
P
Q
R
S
T
U
V
W
X
Y
Z
#misc abbreviations
AB
G
VG
dvs
etc
from
iaf
jfr
kl
kr
mao
mfl
mm
osv
pga
tex
tom
vs

#unified abbreviation list
Acad
Adj
Adm
Adv
Affl
Apr
Art
Asst
Av
Avg
B.ches-du-Rh
Bart
Bco
Bldg
Brig
Bros
C.a
C.p.c.n
Ca
Capt
Cdt
Cf
Ch.-Mme
Chap
Cie
Cmdr
Col
Comdr
Con
Corp
Cpl
DR
DRA
Da
Dec
Dep
Dn
Dr
Dra
Dras
Drs
Eng
Enga
Engas
Engos
Ens
Ets
Euro
Ev
Ex
Excmo
Exmo
Exo
Fa
Fco
Feb
Fig
Fr
Gar
Gen
Gir
Gl
Gov
Hno
Hon
Hosp
Hr
Ilmo
Insp
J.-C
Jan
Jeu
Jr
Jul
Jun
Lda
Lieut
Lt
Lun
MM
MR
MRS
MS
MSc
Maj
Mar
Me
Mej
Mer
Mes
Messrs
Mgr
Mgrs
Mll
Mlle
Mlle(s)
Mme
Mme(s)
Mr
Mrs
Ms
Msgr
Mw
Nov
Npr
Nr
O.d.J
Okt
Op
Ord
Oz
P 
P.D
P.ej
P.p.c
Pas
Pfc
Ph
Prim
Prof
Pte
Pts
Pvt
Rep
Reps
Res
Rev
Revd
Rh
Riv
Rt
S.Em
S.Exc
S.a.r.l
Sen
Sens
Sep
Sept
Sfc
Sgt
SGT
Sl
Sr
Sra
Sras
Srs
Srta
St
ST
Sta
Ste
Sto
Supt
Surg
Tj
Tr
Ud
Uds
V.Exc
Vd
Vda
Vds
Vz
Z.D
Z.D.H
Z.E
Z.Em
Z.H
Z.K.H
Z.K.M
Z.M
a
a./s
a.C
a.g.v
a.l
abrev
abs
ac
acc
acron
adj
adm
adr
adv
alt
anal
anat
angl
appos
apr
apr 
asc
atm
auj
aux
av
avg
avr
b
b.a.o
b.a.p
b.a.r
bacc
bat
bc
bd
bde
bgen
bijv
bijz
br
bv
c 
c.-a-d
c.a.f
c.i
cc
cf
cft
ch
ch.-l
chbre
chbs
chf
col
coll
cpl
cpt
cpte
cta
d
d.c
d.w.z
dcha
dec
def
dem
dep
dept
dhr
dipl
dispo
div
dpto
dr
dr.h.c
dra
dras
drs
ds
dz
e.c
e.g
e.g
e.k
eccles
ecol
econ
ed
ej
env
ep
eq
et
etc
ev
ex
exmo
exo
exp
expo
f.a.c
fa
fam
fasc
fbg
feb
fem
fevr
ff
fl
fol 
fr
fs 
fut
gd
gde
gdes
gds
gen
gl 
grd
h.-t
hab
i.e
i.p.v
i.s.m
i.t.t
i.v.m
ibid
id
imp
ing
ir
iron
itd
itn
itp 
izq
j
janv
jhr
jkvr
jr
l
lat
lex
lgen
lib
lieut
liv
lkol
loc
lof 
m
m.a.w
m.b.t
m.b.v
m.h.o
m.i
m.i.v
maj
mar
mas
max
med
mevr
min
mll
mr
ms
mtr
mtrs 
n
n 
n.f
n.f.pl
n.m
n.m.pl
npr
o
o.b.s
obs
oct
okt
ord 
oz
p
p 
p.a
p.ej
p.ex
p.g.c.d
p.i
p.j
p.m
p.o
p.p
p.p.c.d
p.p.c.m
p.pa
p.pr
pl
plv
poe
pp
pp 
pr
pr 
pres
prev
prof
px
q.s
qqch
qqf
qqn
qqns
r.-de-ch
r.p.m
rc 
rd 
ref
refl
reg
rev
ro 
rte
s
s 
s.a
s.b.f
s.d
s.e 
s.l
s.l.n.d
s.l.p
s.t.p
s.v.p
s/c
sc
sf
sgt
sl
sr
sra
sras
srs
ss 
sto
t
t.s.v.p
tec
tel
terr
tg
tint
tit 
tj
tr
travx
v
v.intr
v.tr
v.w.t
var
vs
vta 
vx
z.v
zool
Št 
št 
